// No Copyright. Vladislav Aleinik, 2020
//=============================================================================
// UART Controller            
//=============================================================================
// - Asyncronously reads instructions from outside
// - Handles all reads from UART buffer
//=============================================================================
// module UartController(
// 	input clk,

// 	input [31:0]local_addr,
// 	input [31:0]write_data
// );

// endmodule