// No Copyright. Vladislav Aleinik, 2020
//=============================================================================
// VGA Controller                 
//=============================================================================
// - Handles All Writes To Video Memory 
// - Asyncronously Renders Video Memory Through VGA 
//=============================================================================
// module VgaController(
// 	input clk,

// 	input [31:0]local_addr,
// 	input [31:0]write_data
// );

// endmodule
